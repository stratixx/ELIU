BJT charakterystyki wej�ciowe

*OPIS UK�ADU 
*tranzystor typu BC547B (NPN) pracujacy w po�aczeniu WE

Q1 2 1 0 BC547B
*    C B E - ko�c�wki tranzystora

V1 1 0 0.5
* �r�d�o napieciowe steruj�ce baz�

V2 2 0 2V
* �r�d�o napi�ciowe na wyj�ciu


* PARAMETRY MODELU TRANZYSTORA NPN 
* 1. linia: parametry materia�owe, statyczne,  i zwi�zane z zale�no�ciami temperaturowymi  
* 2. linia: wzmocnienia pr�dowe, napi�cia Early'ego i wysoki poziom wstrzykiwania
* 3. i 4. rezystancje obszr�w, parametry dynamiczne
  
.model BC547B NPN(Eg=1.11 Is=7.049f Xti=3 Ise=68f Ne=1.576 Isc=12.4f Nc=1.835
+ Bf=400 Br=1 Xtb=1.5 Vaf=62.79 Ikf=81.57m Ikr=3.924 Nk=.4767 
+ Rc=.9747 Cjc=5.25p Mjc=.3147 Vjc=.5697 Fc=.5 
+ Cje=11.5p Mje=.6715 Vje=.5 Tr=10n Tf=410.2p Itf=1.491 Xtf=40.06 Vtf=10)

*Wyznaczenie punktu pracy
.OP

*Analiza DC dla zmiennej warto�ci napi�c UBE przy kilku wartosciach UCE pradu 
.DC LIN  V1 0.5 0.75 0.01  V2 1 10 4


*Zapis do zbioru wyjsciowego
.print DC IC(Q1) IB(Q1) IE(Q1) VB(Q1)

.PROBE
.END
