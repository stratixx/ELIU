BJT cz�stotliwo�ci graniczne

*OPIS UK�ADU 
*tranzystor typu BC547B (NPN) pracujacy w po�aczeniu WE

Q1 2 1 0 BC547B
*    C B E - ko�c�wki tranzystora

I1 0 1 10u
IG 1 0 AC 1u
* �r�d�o pr�dowe zasilaj�ce baz�

V2 2 0 6
* �r�d�o napi�ciowe na wyj�ciu

* PARAMETRY MODELU TRANZYSTORA NPN 
* 1. linia: parametry materia�owe, statyczne,  i zwi�zane z zale�no�ciami temperaturowymi  
* 2. linia: wzmocnienia pr�dowe, napi�cia Early'ego i wysoki poziom wstrzykiwania
* 3. i 4. rezystancje obszr�w, parametry dynamiczne

.model BC547B NPN(Eg=1.11 IS=7.049f Xti=3 Ise=68f Ne=1.576 Isc=12.4f Nc=1.835
+ BF=280 BR=1 Xtb=1.5  Ikf=81.57m Ikr=3.924 Nk=.4767 
+ Rc=.9747 Cjc=5.25p Mjc=.3147 Vjc=.5697 Fc=.5 
+ Cje=11.5p Mje=.6715 Vje=.5 TR=10n TF=420p Itf=1.491 Xtf=40.06 Vtf=10)

*definicja analizy cz�stotliwo�ciowej
.AC DEC 10 10 300meg 

.PRINT AC IC(Q1) IB(Q1)

.OP

.OPTIONS NOPAGE
.PROBE
.END
