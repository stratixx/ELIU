D charakterystyka w przewodzeniu
.WIDTH IN=80 OUT=80

*opis uk�adu: �r�d�o sta�onapi�ciowe oraz dioda p�przewodnikowa
V1 1 0 0.7
D1 1 0 dELIU

*parametry modelu diody
*IS - pr�d nasycenia
*N - wsp�czynnik emisji
*RS - rezystancja szeregowa
*BV - napi�cie przebicia lawinowego
*IBV - pr�d przebicia lawinowego
*CJO -  pojemno�c z��cza przy zerowej polaryzacji
*M - wsp. zale�ny od typy z��cza (z�. skokowe =0.5, liniowe =0.33)
*VJ - potencja� dyfuzyjny z��cza pn
*TT - czas przelotu

.MODEL dELIU D IS=8E-15 RS=1e-10 N=1 BV=10  IBV=1.0E-5  CJO=3P M=0.5 VJ=0.7 TT=0.5N

*definicja analizy sta�onapieciowej oraz zmian RS
.DC V1 0.0001 0.85 0.01 LIN D dELIU(RS) 1e-10 1 0.3

*Zapis do zbioru wyjsciowego
.print DC I(D1)

*punkt pracy
.OP

.OPTIONS NOPAGE
.PROBE
.END
